`ifndef COM
`define COM

class router_common;
  
  static int num_matches = 0;
  static int num_mismatches = 0;
  static int num_packets = 5;
  
endclass

`endif

